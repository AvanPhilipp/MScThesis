----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10/15/2019 12:57:37 PM
-- Design Name: 
-- Module Name: timing_State_Machine - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity timing_State_Machine is
    Port (
    clk: in std_logic;
    rst: in std_logic;
    video_in: in std_logic_vector (7 downto 0);
    video_out: out  std_logic_vector (7 downto 0);
    h_blank: out std_logic;
    v_blank: out std_logic);
end timing_State_Machine;

architecture Behavioral of timing_State_Machine is

type state_type is (vid, v_b, h_b, hv_b);

subtype word16 is std_logic_vector (7 downto 0);
type sh_reg is array (4 downto 0) of word16;

signal v_in_sig: word16;
signal v_out_sig: word16;
signal h_b_reg, v_b_reg: std_logic;
signal shift_reg: sh_reg;
signal state, next_state: state_type;
signal sav_detect: std_logic_vector(3 downto 0);
--signal eav_v_detect: std_logic_vector(4 downto 0);
signal AV_detect: boolean;


begin

v_in_sig<= video_in;
   
Watcher: process (clk)
begin
    if clk'event and clk='1' then
    
        if (rst = '1') then
            state <= vid;
        else
            state <= next_state;
            if(state = vid) then
                video_out <= shift_reg(4);
            else
                video_out <= (others => '0');
            end if;
            h_blank <= h_b_reg;
            v_blank <= v_b_reg;
        end if;
        
--        for i in 0 to 4-2 loop
--            shift_reg(i+1) <= shift_reg(i);
--        end loop;
--        shift_reg(0) <= v_in_sig;
        shift_reg <= shift_reg(shift_reg'left-1 downto 0) & v_in_sig;
     if AV_detect and (shift_reg(0) = x"80" or shift_reg(0) = x"C7") then
        sav_detect(0) <= '1';
    else
        sav_detect(0) <= '0';
    end if;
    sav_detect(sav_detect'left downto 1) <= sav_detect(sav_detect'left-1 downto 0);
--     if AV_detect and (shift_reg(0) = x"B6" or shift_reg(0) = x"F1") then
--        eav_v_detect(0) <= '1';
--    else
--        eav_v_detect(0) <= '0';
--    end if;
--    eav_v_detect(eav_v_detect'left downto 1) <= eav_v_detect(eav_v_detect'left-1 downto 0);
   end if;
end process;

output_decode: process (clk, v_in_sig)
begin
    if state = vid then
        v_out_sig <= v_in_sig;
        h_b_reg <= '0';
        v_b_reg <= '0';
    end if;
    
    if state = v_b then
        v_out_sig <= (others=>'0');
        h_b_reg <= '0';
        v_b_reg <= '1';
    end if;
    if state = h_b then
        v_out_sig <= (others=>'0');
        h_b_reg <= '1';
        v_b_reg <= '0';
    end if;
    if state = hv_b then
        v_out_sig <= (others=>'0');
        h_b_reg <= '1';
        v_b_reg <= '1';
    end if;
end process;


AV_detect <= shift_reg(3)=x"FF" and shift_reg(2)=x"00" and shift_reg(1)=x"00";



next_state_decode: process (shift_reg, sav_detect, AV_detect)
begin
    next_state <= state;
    case (state) is
        when vid =>
            if AV_detect and (shift_reg(0) = x"9D" or shift_reg(0) = x"DA") then
                next_state <= h_b;
            elsif AV_detect and (shift_reg(0) = x"B6" or shift_reg(0) = x"F1")  then
                next_state <= v_b;
            end if;
        when v_b => 
--            if AV_detect and (shift_reg(0) = x"B6" or shift_reg(0) = x"F1") then
--                next_state <= hv_b;
--            elsif shift_reg = x"FF0000AB" or shift_reg = x"FF0000EC"  then
--                next_state <= v_b;

            if sav_detect(3) = '1' then
                next_state <= vid;
            end if;
        when h_b => 
            if sav_detect(3) = '1' then
                next_state <= vid;
--            elsif eav_v_detect(3) = '1' then
--                next_state <= v_b;
            end if;
--        when hv_b => 
--            if AV_detect and (shift_reg(0) = x"80" or shift_reg(0) = x"C7") then
--                next_state <= vid;
--            elsif AV_detect and (shift_reg(0) = x"AB" or shift_reg(0) = x"EC") then
--                next_state <= v_b;
--            end if;
        when others =>
    end case;
end process;




end Behavioral;

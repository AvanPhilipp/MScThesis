----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10/15/2019 03:51:27 PM
-- Design Name: 
-- Module Name: timing_state_machine - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity timing_state_machine is
    Port (
    clk: in std_logic;
    rst: in std_logic;
    video_in: in std_logic_vector (7 downto 0);
    video_out: out  std_logic_vector (7 downto 0);
    h_blank: in std_logic;
    v_blank: in std_logic);
end timing_state_machine;

architecture Behavioral of timing_state_machine is

type state_type is (send_sav, send_h_eav, send_v_eav, blank, video);

subtype word16 is std_logic_vector (7 downto 0);

--type sh_reg_type is array (5 downto 0) of std_logic_vector (7 downto 0);
type sh_reg_type is array (integer range<>) of std_logic_vector (7 downto 0);
type AV_mem_type is array (0 to 15) of word16;

signal state_reg, state_reg_old: state_type:=blank;
signal v_in_sig, v_out_sig: word16;
signal shift_reg: sh_reg_type(5 downto 0);
signal h_b_reg, h_b_reg_old, v_b_reg, v_b_reg_old : std_logic;
signal blank_count: std_logic_vector (4 downto 0);
signal sav_counter: unsigned (1 downto 0);
signal eav_counter: unsigned (3 downto 0);

signal AV_memory: AV_mem_type := (  x"FF",x"00", x"00",x"80",
                                    x"FF",x"00", x"00",x"9D",
                                    x"FF",x"00", x"00",x"AB",
                                    x"FF",x"00", x"00",x"B6");
signal AV_memory_reg: word16;
signal AV_memory_reg_shifted: sh_reg_type (3 downto 0);


begin

Watcher: process (clk) begin
    if clk'event and clk='1' then
        
        --Incoming signal to register
        v_in_sig <= video_in;
        h_b_reg <= h_blank;
        v_b_reg <= v_blank;
        state_reg_old <= state_reg;
        
        --Decode Output
        if state_reg_old = blank then
--            video_out <= (others => '0');
            video_out <=  shift_reg(shift_reg'left);
        elsif state_reg_old = send_sav then
             video_out <= AV_memory_reg;
       elsif state_reg = send_h_eav or state_reg = send_v_eav then
            if eav_counter(3 downto 2) = "00" or eav_counter = 4 then
                video_out <=  shift_reg(shift_reg'left);
            else
                video_out <= AV_memory_reg;
            end if;
--            video_out <= AV_memory_reg;
--            shift_reg(shift_reg'left) <= AV_memory_reg;
        elsif state_reg_old = video then
            video_out <= shift_reg(shift_reg'left);
        else
            video_out <= (others => '0');
        end if;
        
        --Shift registers
        shift_reg <= shift_reg(shift_reg'left-1 downto 0) & v_in_sig;
        AV_memory_reg_shifted <= AV_memory_reg_shifted(AV_memory_reg_shifted'left-1 downto 0) & AV_memory_reg;
        
        -- Blanking signal detect
        h_b_reg_old <= h_b_reg;
        v_b_reg_old <= v_b_reg;
        
        -- Next State Logic
        case (state_reg) is
            when blank =>
                if h_b_reg_old = '1' and h_b_reg = '0' and v_b_reg = '0' then
                    state_reg <= send_sav;
                end if;
            when send_sav =>
                if sav_counter = 3 then
                    state_reg <= video;
                end if;
            when video =>
                if h_b_reg_old = '0' and h_b_reg = '1' then
                    if v_b_reg = '1' then
                        state_reg <= send_v_eav;
                    else
                        state_reg <= send_h_eav;
                    end if;
                end if;
            when send_v_eav | send_h_eav =>
                if eav_counter = 8 then
                    state_reg <= blank;
                end if;
            when others =>
                state_reg <= blank;
        end case;
            
            
        -- Active Video Counter
        if state_reg = send_sav then 
            sav_counter <= sav_counter + 1;
        else
            sav_counter <= (others => '0');
        end if;
        
        if state_reg = send_v_eav or state_reg = send_h_eav then
            eav_counter <= eav_counter + 1;
        else
            eav_counter <= (others => '0');
        end if;
        
        
        --Memory Adderss Decode
        if state_reg = send_sav then
            AV_memory_reg <= AV_memory(to_integer("00" & sav_counter));
        elsif state_reg = send_h_eav then 
            AV_memory_reg <= AV_memory(to_integer("01" & eav_counter(1 downto 0)));
        elsif state_reg = send_v_eav then 
            AV_memory_reg <= AV_memory(to_integer("10" & eav_counter(1 downto 0)));
        end if;
        
--        --Memory Adderss Decode
--        if state_reg = send_sav then
--            AV_memory_reg <= AV_memory(to_integer("00" & av_counter));
--        elsif h_b_reg = '1' then 
--            AV_memory_reg <= AV_memory(to_integer("01" & av_counter));
--        elsif h_b_reg_old = '0' and h_b_reg = '1' and v_b_reg = '1' then
--            AV_memory_reg <= AV_memory(to_integer("10" & av_counter));
--        end if;

   end if;
end process;


end Behavioral;


